module and_8_entradas(e,z);

input [7:0] e;

output z;

and (z,e[0],e[1],e[2],e[3],e[4],e[5],e[6],e[6],e[7]);

endmodule 

module estagio_ula_1000(ack_in);

input ack_in;

estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();
estagio_ula();

endmodule 
